// Code your testbench here
// or browse Examples
module array;
  int arr[3][5][5]='{'{'{1,2,3,4,5},
                   '{10,20,30,40,50},
                   '{12,22,53,49,45},
                   '{85,34,66,2,0},
                     '{2,3,4,5,6}},
                    '{'{1,2,3,4,5},
                   '{10,20,30,40,50},
                   '{12,22,53,49,45},
                   '{85,34,66,2,0},
                      '{2,3,4,5,6}},
  				        	'{'{1,2,3,4,5},
                   '{10,20,30,40,50},
                   '{12,22,53,49,45},
                   '{85,34,66,2,0},
                      '{2,3,4,5,6}}};
  			
  initial begin
    foreach(arr[i,j,k])begin
      $display("array[%0d][%0d][%0d]=%0d",i,j,k,arr[i][j][k]);
   end
  end
endmodule
