class A;
  int a;
  int i;
  mailbox m;
  
  function new(mailbox m1);
  this.m = m1;
  endfunction
  
  task check();
    if(m==null)
      $display("Mailbox is not full");
    else
      $display("Mailbox is created");
    
    for(i=0;i<3;i++)begin
    a++;
      m.put(a);
      $display("value of a = %0d",a);
    end
  endtask
endclass

module tb;
  A a1;
  mailbox main = new(3);
  initial begin
    a1 = new(main);
    a1.check();
  end
endmodule
/*Mailbox is created
value of a = 1
value of a = 2
value of a = 3*/
